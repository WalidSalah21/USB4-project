`timescale 1ns/1ps

module  pulse_sync_3bit_tb ;

/////////////////////////////////////////////////////////
///////////////////// Parameters ////////////////////////
/////////////////////////////////////////////////////////

parameter Clock_PERIOD_a = 10 ; //fast clock
parameter Clock_PERIOD_b = 10000 ; //slow clock


/////////////////////////////////////////////////////////
//////////////////// DUT Signals ////////////////////////
/////////////////////////////////////////////////////////

reg        clk_a_tb;
reg        clk_b_tb;
reg        rst_tb;
reg  [2:0] sig_4bit_tb;
wire       busy_tb;
wire [2:0] sig_sync_4bit_tb;


////////////////////////////////////////////////////////
////////////////// initial block /////////////////////// 
////////////////////////////////////////////////////////

initial 
 begin
 
 // t=0
clk_a_tb = 0;
clk_b_tb = 0;
rst_tb = 0;
sig_4bit_tb = 'h0;

#(Clock_PERIOD_a) 
rst_tb = 1;

@ (posedge clk_a_tb)
sig_4bit_tb = 'h6;

@ (posedge clk_a_tb)
sig_4bit_tb = 'h0;

 end


////////////////////////////////////////////////////////
////////////////// Clock Generator  ////////////////////
////////////////////////////////////////////////////////

always #(Clock_PERIOD_a/2)  clk_a_tb = ~clk_a_tb ;
always #(Clock_PERIOD_b/2)  clk_b_tb = ~clk_b_tb ;


////////////////////////////////////////////////////////
/////////////////// DUT Instantation ///////////////////
////////////////////////////////////////////////////////

pulse_sync_3bit DUT
(
.sig_3bit(sig_4bit_tb), 
.rst(rst_tb), 
.clk_a(clk_a_tb), 
.clk_b(clk_b_tb), 
.sig_sync_3bit(sig_sync_4bit_tb),
.busy(busy_tb)
);

endmodule