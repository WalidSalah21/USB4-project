package top_elec;

`include "path_to_your_file/elec_layer_tr.sv";
`include "elec_layer_generator.sv";
`include "elec_layer_driver.sv";
`include "elec_layer_monitor.sv";

endpackage: top_elec